library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.CONV_STD_LOGIC_VECTOR;
use work.HermesPackage.all;

entity topNoC is
end;

architecture topNoC of topNoC is

	signal clock : regNrot;
	signal reset, finish : std_logic;
	signal clock_rx, rx, credit_o: regNrot;
	signal clock_tx, tx, credit_i: regNrot;
	signal data_in, data_out : arrayNrot_regflit;

	signal address1, data1 : std_logic_vector(15 downto 0);
	signal ce1 : std_logic;

	constant pck1 : service_request_packet := (
		x"C122", x"0003", service_request, x"0000", x"000A"
	);
	-- C122 (C = peripheral communication; 1 = north port; 22 = target PE coord)
	-- 0003 = number of flits
	-- 1001 = request service
	-- 0000 = (first part is reserved, second part 00 = source PE)
	-- 000A = task id

	constant pck2 : service_request_packet := (
		x"C122", x"0003", x"1001", x"0000", x"000B"
	);

begin
	reset <= '1', '0' after 15 ns;

	-- clock process of router N0000
	process
	begin
		clock(N0000) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0100
	process
	begin
		clock(N0100) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0200
	process
	begin
		clock(N0200) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0001
	process
	begin
		clock(N0001) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0101
	process
	begin
		clock(N0101) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0201
	process
	begin
		clock(N0201) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0002
	process
	begin
		clock(N0002) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0102
	process
	begin
		clock(N0102) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	-- clock process of router N0202
	process
	begin
		clock(N0202) <= '1', '0' after 10 ns;
		wait for 20 ns;
	end process;

	NOC: Entity work.NOC
	port map(
		clock         => clock,
		reset         => reset,
		clock_rxLocal => clock_rx,
		rxLocal       => rx,
		data_inLocal  => data_in,
		credit_oLocal => credit_o,
		clock_txLocal => clock_tx,
		txLocal       => tx,
		data_outLocal => data_out,
		credit_iLocal => credit_i);

	--com00: Entity work.outmodule
	--port map(
	--	clock       => clock(N0000),
	--	reset       => reset,
	--	finish      => finish,
	--	inClock0    => clock_tx(N0000),
	--	inTx0       => tx(N0000),
	--	inData0     => data_out(N0000),
	--	outCredit0  => credit_i(N0000),
	--	inClock1    => clock_tx(N0100),
	--	inTx1       => tx(N0100),
	--	inData1     => data_out(N0100),
	--	outCredit1  => credit_i(N0100),
	--	inClock2    => clock_tx(N0200),
	--	inTx2       => tx(N0200),
	--	inData2     => data_out(N0200),
	--	outCredit2  => credit_i(N0200),
	--	inClock3    => clock_tx(N0001),
	--	inTx3       => tx(N0001),
	--	inData3     => data_out(N0001),
	--	outCredit3  => credit_i(N0001),
	--	inClock4    => clock_tx(N0101),
	--	inTx4       => tx(N0101),
	--	inData4     => data_out(N0101),
	--	outCredit4  => credit_i(N0101),
	--	inClock5    => clock_tx(N0201),
	--	inTx5       => tx(N0201),
	--	inData5     => data_out(N0201),
	--	outCredit5  => credit_i(N0201),
	--	inClock6    => clock_tx(N0002),
	--	inTx6       => tx(N0002),
	--	inData6     => data_out(N0002),
	--	outCredit6  => credit_i(N0002),
	--	inClock7    => clock_tx(N0102),
	--	inTx7       => tx(N0102),
	--	inData7     => data_out(N0102),
	--	outCredit7  => credit_i(N0102),
	--	inClock8    => clock_tx(N0202),
	--	inTx8       => tx(N0202),
	--	inData8     => data_out(N0202),
	--	outCredit8  => credit_i(N0202));

	clock_rx(N0100) <= '0';
	rx(N0100) <= '0';
	
	clock_rx(N0200) <= '0';
	rx(N0200) <= '0';
	
	clock_rx(N0001) <= '0';
	rx(N0001) <= '0';
	
	clock_rx(N0101) <= '0';
	rx(N0101) <= '0';
	
	clock_rx(N0201) <= '0';
	rx(N0201) <= '0';
	
	clock_rx(N0002) <= '0';
	rx(N0002) <= '0';
	
	clock_rx(N0102) <= '0';
	rx(N0102) <= '0';
	
	clock_rx(N0202) <= '0';
	rx(N0202) <= '0';


	clock_rx(N0000) <= clock(N0000); --clock to inject data -the same of the router

	process(reset, clock(N0000))
	begin
		if reset = '1' then
			rx(N0000) <= '0';
		elsif clock(N0000)'event and clock(N0000)='1' then
			if ce1 = '1' and address1 = x"FFFF" then
				rx(N0000) <= '1';
				data_in(N0000) <= data1;
			elsif credit_o(N0000) = '1' then --important: flow control
				rx(N0000) <= '0';
			end if;
		end if;
	end process;

	address1 <= x"FFFF"; --address generated by the processor

	process
		variable i : integer:= 0;
	begin
		ce1 <= '0';
		wait for 500 ns; --time between packets
		i := 0;

		while i < 5 loop
			if credit_o(N0000)='1' then --important: flow control
				data1 <= pck1(i); --simulate a write( pck(i), address_noc)
				ce1  <= '1';
				wait for 20 ns;
				ce1  <= '0';
				wait for 20 ns;
				i := i + 1;
			else
				wait for 20 ns;
			end if;
		end loop;

		wait for 500 ns; --time between packets
		i := 0;
		while i < 5 loop
			if credit_o(N0000)='1' then --important: flow control
				data1 <= pck2(i); --simulate a write( pck(i), address_noc)
				ce1  <= '1';
				wait for 20 ns;
				ce1  <= '0';
				wait for 20 ns;
				i := i + 1;
			else
				wait for 20 ns;
			end if;
		end loop;

		wait for 2000 ns; --time between packets
	end process;

end topNoC;
